module helloworld;

initial begin
	$display ("helloworld!!\n");
	#10 $finish;
end
endmodule

